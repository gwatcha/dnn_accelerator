module tb_wordcopy();
endmodule: tb_wordcopy
