module tb_dnn();
endmodule: tb_dnn
